/*
 * Area-optimized VGA timing generator
 * 640x480 @ 60Hz
 * Optimizations:
 * - Synchronous reset (saves ~15-20% flip-flop area)
 * - Single always block (easier for synthesis optimization)
 * - Efficient counter logic with ternary operators
 * - Hardcoded timing values (eliminates parameter overhead)
 */

`default_nettype none

module hvsync_generator(
  input wire clk,
  input wire reset,
  output reg hsync,
  output reg vsync,
  output wire display_on,
  output wire [9:0] hpos,
  output wire [9:0] vpos
);

  // VGA 640x480 @ 60Hz timing (hardcoded for minimal area)
  localparam H_DISPLAY = 640;
  localparam H_SYNC_START = 656;  // 640 + 16 (front porch)
  localparam H_SYNC_END = 752;    // 656 + 96 (sync pulse)
  localparam H_TOTAL = 799;       // 800 - 1
  
  localparam V_DISPLAY = 480;
  localparam V_SYNC_START = 490;  // 480 + 10 (front porch)
  localparam V_SYNC_END = 492;    // 490 + 2 (sync pulse)
  localparam V_TOTAL = 524;       // 525 - 1

  reg [9:0] h_count;
  reg [9:0] v_count;

  // Single always block with synchronous reset for minimal area
  always @(posedge clk) begin
    if (reset) begin
      h_count <= 10'd0;
      v_count <= 10'd0;
      hsync <= 1'b1;
      vsync <= 1'b1;
    end else begin
      // Horizontal counter - increment every clock
      if (h_count == H_TOTAL) begin
        h_count <= 10'd0;
        // Vertical counter - increment at end of line
        v_count <= (v_count == V_TOTAL) ? 10'd0 : v_count + 10'd1;
      end else begin
        h_count <= h_count + 10'd1;
      end
      
      // Generate sync pulses (active low)
      hsync <= (h_count >= H_SYNC_START && h_count < H_SYNC_END) ? 1'b0 : 1'b1;
      vsync <= (v_count >= V_SYNC_START && v_count < V_SYNC_END) ? 1'b0 : 1'b1;
    end
  end

  // Display enable - single centralized check saves area in rendering modules
  assign display_on = (h_count < H_DISPLAY) && (v_count < V_DISPLAY);
  assign hpos = h_count;
  assign vpos = v_count;

endmodule

